package hippo_decoder_ConfigPkg;

    // CSR Related
    typedef logic [12-1:0] CsrAddr;

endpackage
//# sourceMappingURL=config_pkg.sv.map
