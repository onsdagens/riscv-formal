`ifdef __veryl_test_hippomenes_veryl_alu__
    `ifdef __veryl_wavedump_hippomenes_veryl_alu__
        module __veryl_wavedump;
            initial begin
                $dumpfile("alu.vcd");
                $dumpvars();
            end
        endmodule
    `endif
`ifndef SYNTHESIS
import hippo_alu_veryl_ALUPackage::*;
module tb_alu;

  logic [31:0] a;
  logic [31:0] b;
  ALUOp op;
  logic sub_arith;

  logic [31:0] res;

  hippo_alu_veryl_HippoALU dut (
      .a(a),
      .b(b),
      .op(op),
      .sub_arith(sub_arith),
      .res(res)
  );

  initial begin
    $dumpfile("alu.fst");
    $dumpvars;

    a = 3;
    b = 5;
    op = ALUOp_ALU_ADD;
    sub_arith = 0;

    #10;
    assert (res == 8) $display("3 + 5 = 8");
    else $error();

    a  = 3;  // 011
    b  = 5;  // 101
    op = ALUOp_ALU_SLT;
    #10;
    assert (res == 1) $display("(3 < 5) -> true");
    else $error();

    a  = -3;
    b  = 5;
    op = ALUOp_ALU_SLT;
    #10;
    assert (res == 1) $display("signed (-3 < 5) -> true");
    else $error();

    a  = -3;
    b  = 5;
    op = ALUOp_ALU_SLTU;
    #10;
    assert (res == 0) $display("unsigned (-3 < 5) -> false");
    else $error();

    a  = -3;
    b  = -5;
    op = ALUOp_ALU_SLT;
    #10;
    assert (res == 0) $display("signed (-3 < -5) -> false");
    else $error();

    a  = -3;
    b  = -5;
    op = ALUOp_ALU_SLTU;
    #10;
    assert (res == 0) $display("unsigned (-3 < -5) -> false");
    else $error();

    a  = 3;
    b  = -5;
    op = ALUOp_ALU_SLTU;
    #10;
    assert (res == 1) $display("unsigned (3 < -5) -> true");
    else $error();

    a  = 3;
    b  = -5;
    op = ALUOp_ALU_SLT;
    #10;
    assert (res == 0) $display("signed (3 < -5) -> false");
    else $error();

    // shifting
    a  = 3;
    b  = 2;
    op = ALUOp_ALU_SLL;
    #10;
    assert (res == 12) $display("(3 << 2) = 12");
    else $error();

    a = 12;
    b = 2;
    op = ALUOp_ALU_SR;
    sub_arith = 0;  // shift right logic
    #10;
    assert (res == 3) $display("unsigned (12 >> 2) = 3");
    else $error();

    a = -12;
    b = 2;
    op = ALUOp_ALU_SR;
    sub_arith = 0;
    #10;
    assert(res == 'h3ffffffd) $display("unsigned (-12 >> 2) = 0x3ffffffd");
    else $error("logical right shift fail");

    a = 12;
    b = 2;
    op = ALUOp_ALU_SR;
    sub_arith = 1;  // shift right arithmetic
    #10;
    assert (res == 3) $display("signed (12 >> 2) = 3");
    else $error();

    a = -12;
    b = 2;
    op = ALUOp_ALU_SR;
    sub_arith = 1;  // shift right arithmetic
    #10;
    //assert (res == -3) $display("signed(-12 >>> 2) = -3");
    //else $error("arithmetic right shift fail res = %h", res);

    #10 $finish;

  end
endmodule
`endif
`endif
//# sourceMappingURL=test_bench.sv.map
