package hippo_alu_veryl_ALUPackage;
    typedef enum logic [3-1:0] {
        ALUOp_ALU_ADD,
        ALUOp_ALU_SLL,
        ALUOp_ALU_SLT,
        ALUOp_ALU_SLTU,
        ALUOp_ALU_XOR,
        ALUOp_ALU_SR,
        ALUOp_ALU_OR,
        ALUOp_ALU_AND
    } ALUOp;
endpackage
//# sourceMappingURL=alu_pkg.sv.map
